library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity memoria is
	port(
		control: in std_logic;
		clock: in std_logic; --SeÃƒÆ’Ã‚Â±al de reloj
		s_22: in std_logic := '1'; --s_22=1 ESCRITURA,s_22=0 LECTURA
		address: in integer range 0 to 65535; --16 direcciones codificadas por 5 bits
		data_in: in std_logic_vector (7 downto 0); --Ancho de palabra de 8 bits
		data_out: out std_logic_vector (7 downto 0)); --Salida de datos
end memoria;

architecture rtl of memoria is
	-- Build a 2-D array type for the RAM
	subtype word_t is std_logic_vector(7 downto 0);
	type datos is array (53759 downto 0) of word_t;
	
	-- Declare the RAM signal.
	signal ram : datos := (
		0 => "01100100",
		1 => "00000001",
		2 => "00000000",
		3 => "00000000",
		4 => "00000000",
		5 => "00000000",
		6 => "00000000",
		7 => "00000000",
		8 => "00000000",
		9 => "00000000",
		10 => "00000000",
		11 => "00000000",
		12 => "00000000",
		13 => "00000000",
		14 => "00000000",
		15 => "00000000",
		16 => "00000000",
		17 => "00000000",
		18 => "00000000",
		19 => "00000000",
		20 => "00000000",
		21 => "00000000",
		22 => "00000000",
		23 => "00000000",
		24 => "00000000",
		25 => "00000000",
		26 => "00000000",
		27 => "00000000",
		28 => "00000000",
		29 => "00000000",
		30 => "00000000",
		31 => "00000000",
		32 => "00000000",
		33 => "00000000",
		34 => "00000000",
		35 => "00000000",
		36 => "00000000",
		37 => "00000000",
		38 => "00000000",
		39 => "00000000",
		40 => "00000000",
		41 => "00000000",
		42 => "00000000",
		43 => "00000000",
		44 => "00000000",
		45 => "00000000",
		46 => "00000000",
		47 => "00000000",
		48 => "00000000",
		49 => "00000000",
		50 => "00000000",
		51 => "00000000",
		52 => "00000000",
		53 => "00000000",
		54 => "00000000",
		55 => "00000000",
		56 => "00000000",
		57 => "00000000",
		58 => "00000000",
		59 => "00000000",
		60 => "00000000",
		61 => "00000000",
		62 => "00000000",
		63 => "00000000",
		64 => "00000000",
		65 => "00000000",
		66 => "00000000",
		67 => "00000000",
		68 => "00000000",
		69 => "00000000",
		70 => "00000000",
		71 => "00000000",
		72 => "00000000",
		73 => "00000000",
		74 => "00000000",
		75 => x"00",
		76 => x"02",
		77 => x"72",
		78 => x"00",
		79 => x"00",
		80 => x"C3",
		81 => x"00",
		82 => x"28",
		83 => x"36",
		84 => x"00",
		85 => x"92",
		86 => x"36",
		87 => x"00",
		88 => x"A8",
		89 => x"43",
		90 => x"28",
		91 => x"00",
		92 => x"63",
		93 => x"36",
		94 => x"00",
		95 => x"B4",
		96 => x"35",
		97 => x"00",
		98 => x"8A",
		99 => x"36",
		100 => x"00",
		101 => x"CA",
		102 => x"36",
		103 => x"00",
		104 => x"FB",
		105 => x"27",
		106 => x"00",
		107 => x"72",
		108 => x"33",
		109 => x"00",
		110 => x"07",
		111 => x"34",
		112 => x"00",
		113 => x"08",
		114 => x"71",
		115 => x"00",
		116 => x"07",
		117 => x"B1",
		118 => x"00",
		119 => x"08",
		120 => x"79",
		121 => x"00",
		122 => x"01",
		123 => x"8B",
		124 => x"00",
		125 => x"18",
		126 => x"00",
		127 => x"86",
		128 => x"15",
		129 => x"00",
		130 => x"63",
		131 => x"35",
		132 => x"00",
		133 => x"8A",
		134 => x"91",
		135 => x"28",
		136 => x"00",
		137 => x"63",
		138 => x"71",
		139 => x"00",
		140 => x"04",
		141 => x"B1",
		142 => x"00",
		143 => x"03",
		144 => x"1F",
		145 => x"10",
		146 => x"31",
		147 => x"00",
		148 => x"03",
		149 => x"31",
		150 => x"00",
		151 => x"04",
		152 => x"31",
		153 => x"00",
		154 => x"05",
		155 => x"31",
		156 => x"00",
		157 => x"06",
		158 => x"31",
		159 => x"00",
		160 => x"02",
		161 => x"31",
		162 => x"00",
		163 => x"07",
		164 => x"31",
		165 => x"00",
		166 => x"08",
		167 => x"37",
		168 => x"41",
		169 => x"01",
		170 => x"72",
		171 => x"00",
		172 => x"06",
		173 => x"71",
		174 => x"00",
		175 => x"00",
		176 => x"72",
		177 => x"00",
		178 => x"04",
		179 => x"37",
		180 => x"41",
		181 => x"F7",
		182 => x"81",
		183 => x"0F",
		184 => x"C1",
		185 => x"08",
		186 => x"72",
		187 => x"00",
		188 => x"03",
		189 => x"B2",
		190 => x"00",
		191 => x"04",
		192 => x"72",
		193 => x"00",
		194 => x"05",
		195 => x"B2",
		196 => x"00",
		197 => x"06",
		198 => x"F2",
		199 => x"00",
		200 => x"02",
		201 => x"37",
		202 => x"71",
		203 => x"00",
		204 => x"03",
		205 => x"B1",
		206 => x"00",
		207 => x"04",
		208 => x"78",
		209 => x"00",
		210 => x"05",
		211 => x"BA",
		212 => x"00",
		213 => x"06",
		214 => x"72",
		215 => x"00",
		216 => x"03",
		217 => x"B2",
		218 => x"00",
		219 => x"04",
		220 => x"FD",
		221 => x"00",
		222 => x"04",
		223 => x"7D",
		224 => x"00",
		225 => x"03",
		226 => x"71",
		227 => x"00",
		228 => x"00",
		229 => x"72",
		230 => x"00",
		231 => x"13",
		232 => x"BF",
		233 => x"00",
		234 => x"03",
		235 => x"B0",
		236 => x"00",
		237 => x"10",
		238 => x"36",
		239 => x"01",
		240 => x"0E",
		241 => x"FF",
		242 => x"00",
		243 => x"16",
		244 => x"F0",
		245 => x"00",
		246 => x"05",
		247 => x"73",
		248 => x"00",
		249 => x"02",
		250 => x"37",
		251 => x"71",
		252 => x"00",
		253 => x"03",
		254 => x"B1",
		255 => x"00",
		256 => x"04",
		257 => x"79",
		258 => x"00",
		259 => x"05",
		260 => x"BB",
		261 => x"00",
		262 => x"06",
		263 => x"72",
		264 => x"00",
		265 => x"07",
		266 => x"B2",
		267 => x"00",
		268 => x"08",
		269 => x"37",
		270 => x"C1",
		271 => x"18",
		272 => x"31",
		273 => x"00",
		274 => x"16",
		275 => x"31",
		276 => x"00",
		277 => x"17",
		278 => x"31",
		279 => x"00",
		280 => x"14",
		281 => x"31",
		282 => x"00",
		283 => x"15",
		284 => x"36",
		285 => x"01",
		286 => x"33",
		287 => x"36",
		288 => x"01",
		289 => x"46",
		290 => x"25",
		291 => x"01",
		292 => x"2E",
		293 => x"73",
		294 => x"00",
		295 => x"16",
		296 => x"72",
		297 => x"00",
		298 => x"14",
		299 => x"B2",
		300 => x"00",
		301 => x"15",
		302 => x"64",
		303 => x"28",
		304 => x"01",
		305 => x"1C",
		306 => x"37",
		307 => x"BE",
		308 => x"00",
		309 => x"12",
		310 => x"7E",
		311 => x"00",
		312 => x"13",
		313 => x"7E",
		314 => x"00",
		315 => x"14",
		316 => x"7E",
		317 => x"00",
		318 => x"15",
		319 => x"BE",
		320 => x"00",
		321 => x"16",
		322 => x"7E",
		323 => x"00",
		324 => x"17",
		325 => x"37",
		326 => x"71",
		327 => x"00",
		328 => x"14",
		329 => x"79",
		330 => x"00",
		331 => x"10",
		332 => x"B1",
		333 => x"00",
		334 => x"15",
		335 => x"BB",
		336 => x"00",
		337 => x"11",
		338 => x"37",

        -- Finalizando a memoria com zeros
        others => "00000000"
    );
	
	--signal posicion:integer;
	-- Register to hold the address
	signal addr_reg : integer range 0 to 63;
begin
	--posicion<= to_integer(unsigned(address));
	process (clock)
	begin
		if(falling_edge(clock)) then
			if(s_22 = '1') then
				if(control = '1') then
					ram(address) <= data_in;
				end if;
			end if;
		end if;
	end process;
	
	data_out <= ram(address);
	
end rtl;