-- Memoria de microcodigo
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity mem_micro_cod is
    port (
        clk : in std_logic;
        addr : in std_logic_vector(7 downto 0);
        data : out std_logic_vector(23 downto 0)
    );
end mem_micro_cod;

architecture rtl of mem_micro_cod is
    type mem_type is array (0 to 255) of std_logic_vector(23 downto 0);
    signal mem : mem_type := (
		0  => "000000011000000000000001",  --- Instrucion de comienzo
        1  => "000000000000000100000001",
        2  => "010000000000000000000011",

        16 => "000000000000000100000001",  --- Direccionamiento Inherente
        17 => "010000000000000000000001",
        18 => "000000101011000000000111",

        32 => "000000000000000100000001",  --- Direccionamiento Inmediato
        33 => "010000000000000000000001",
        34 => "000000101000000000000001",
        35 => "000000000000000100000001",
        36 => "000000101000000000000111",

        48 => "000000000000000100000001",  --- Direccionamiento Directo
        49 => "010000000000000000000001",
        50 => "000000101000000000000001",
        51 => "000000000000000100000001",
        52 => "000010000000000000000001",
        53 => "000000101000000000000001",
        54 => "000000000000000100000001",
        55 => "000001000000010000000001",
        56 => "000000000000010100000001",
        57 => "000000101000000011000111",

        64 => "000000000000000100000001",  --- Direccionamiento Indexado
        65 => "010000000000000000000001",
        66 => "000000101000000000000001",
        67 => "000000000000000100000001",
        68 => "101000000000000000000001",
        69 => "001000101000000000000001",
        70 => "001000000000000100000001",
        71 => "001100000000000000000001",
        72 => "001000000000100100000001",
        73 => "001000101000000011000111",

        80 => "000000000000000100000001",  --- Instruccion de Salto
        81 => "010000000000000000000001",
        82 => "000000101000000000000001",
        83 => "000000000000000100000001",
        84 => "000010000000000000000001",
        85 => "000000101000000000000001",
        86 => "000000000000000100000001",
        87 => "000001000000010000000001",
        88 => "000000111100000000000011",
        
        96 => "000000000000000100000001",  --- Instruccion de Subrutina
        97 => "010000000000000000000001",
        98 => "000000101000000000000001",
        99 => "000000000000000100000001",
        100 => "000010000000000000000001",
        101 => "000000101000000000000001",
        102 => "000000000000000100000001",
        103 => "000001000000010000000001",
        104 => "000000101000000000000001",
        105 => "000000000001000000000001",
        106 => "000000000000110100000001",
        107 => "000000000000000010110001",
        108 => "000000000001000000000001",
        109 => "000000000000110100000001",
        110 => "000000000000000010111001",
        111 => "000000011100000000000011",

        112 => "000000000000000100000001",  --- Instruccion de Retorno de Subrutina
        113 => "010000000000000000000001",
        114 => "000000000000110100000001",
        115 => "000001000000000000000001",
        116 => "000000000001000000000001",
        117 => "000000000000110100000001",
        118 => "000010000000000000000001",
        119 => "000000000001000000000001",
        120 => "000000011100000000000011",

        128 => "000000000000000100000001",  --- Instruccion de Guardado de punteros
        129 => "010000000000000000000001",
        130 => "000000101000000000000001",
        131 => "000000000000000100000001",
        132 => "000010000000000000000001",
        133 => "000000101000000000000001",
        134 => "000000000000000100000001",
        135 => "000001000000000000000001",
        136 => "000000000000010100000001",
        137 => "000000000000000011110001",
        138 => "000000000000001000000001",
        139 => "000000000000000011111001",
        140 => "000000101000000000000011",

        144 => "000000000000000100000001",  --- Instruccion de Carga de punteros Inmediata
        145 => "010000000000000000000001",
        146 => "000000101000000000000001",
        147 => "000000000000000100000001",
        148 => "000010000000000000000001",
        149 => "000000101000000000000001",
        150 => "000000000000000100000001",
        151 => "000001000000000000000001",
        152 => "000000101011000000000011",

        160 => "000000000000000100000001",  --- Instruccion de Carga de punteros Directa
        161 => "010000000000000000000001",
        162 => "000000101000000000000001",
        163 => "000000000000000100000001",
        164 => "000010000000000000000001",
        165 => "000000101000000000000001",
        166 => "000000000000000100000001",
        167 => "000001000000000000000001",
        168 => "000000000000010100000001",
        169 => "000010000000000000000001",
        170 => "000000000000001000000001",
        171 => "000001000000000000000001",
        172 => "000000101011000000000011",

        176 => "000000000000000100000001",  --- Instruccion de Guardado en pila de Acumulador
        177 => "010000000000000000000001",
        178 => "000000000001000000000001",
        179 => "000000000000110100000001",
        180 => "000000101000000011001111",

        192 => "000000000000000100000001",  --- Instruccion de Guardado en pila de Punteros
        193 => "010000000000000000000001",
        194 => "000000000001000000000001",
        195 => "000000000000110100000001",
        196 => "000000000000000010010001",
        197 => "000000000001000000000001",
        198 => "000000000000110100000001",
        199 => "000000000000000010011001",
        200 => "000000101000000000000011",

        208 => "000000000000000100000001",  --- Instruccion de Recuperado de pila Acumulador
        209 => "010000000000000000000001",
        210 => "000000000000110100000001",
        211 => "000000101001000000000111",

        224 => "000000000000000100000001",  --- Instruccion de Recuperado de pila Punteros
        225 => "010000000000000000000001",
        226 => "000000000000110100000001",
        227 => "000001000000000000000001",
        228 => "000000000001000000000001",
        229 => "000000000000110100000001",
        230 => "000010000000000000000001",
        231 => "000000101010000000000001",
        232 => "000000000001000000000011",

        -- Finalizando a memoria com zeros
        others => "000000000000000000000001"
    );

begin
    process(clk)
    begin
        if rising_edge(clk) then
            data <= mem(to_integer(unsigned(addr)));
        end if;
    end process;
end rtl;