-- Memoria de microcodigo
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity mem_micro_cod is
    port (
        clk : in std_logic;
        addr : in std_logic_vector(7 downto 0);
        data : out std_logic_vector(24 downto 0)
    );
end mem_micro_cod;

architecture rtl of mem_micro_cod is
    type mem_type is array (0 to 255) of std_logic_vector(24 downto 0);
    signal mem : mem_type := (
		0  => "0000000011000000000000001",  --- Instrucion de comienzo
        1  => "0000000000000000100000001",
        2  => "0010000000000000000000011",

        16 => "0000000000000000100000001",  --- Direccionamiento Inherente
        17 => "0010000000000000000000001",
        18 => "0000000101011000000000111",

        32 => "0000000000000000100000001",  --- Direccionamiento Inmediato
        33 => "0010000000000000000000001",
        34 => "0000000101000000000000001",
        35 => "0000000000000000100000001",
        36 => "0000000101000000000000111",

        48 => "0000000000000000100000001",  --- Direccionamiento Directo
        49 => "0010000000000000000000001",
        50 => "0000000101000000000000001",
        51 => "0000000000000000100000001",
        52 => "0000010000000000000000001",
        53 => "0000000101000000000000001",
        54 => "0000000000000000100000001",
        55 => "0000001000000010000000001",
        56 => "0000000000000010100000001",
        57 => "0000000101000000011000111",

        64 => "0000000000000000100000001",  --- Direccionamiento Indexado
        65 => "0010000000000000000000001",
        66 => "0000000101000000000000001",
        67 => "0000000000000000100000001",
        68 => "0100000000000000000000001",
        69 => "0001000101000000000000001",
        70 => "0001000000000000100000001",
        71 => "0001100000000000000000001",
        72 => "0001000000000100100000001",
        73 => "0001000101000000011000111",

        80 => "0000000000000000100000001",  --- Instruccion de Salto
        81 => "0010000000000000000000001",
        82 => "0000000101000000000000001",
        83 => "0000000000000000100000001",
        84 => "0000010000000000000000001",
        85 => "0000000101000000000000001",
        86 => "0000000000000000100000001",
        87 => "0000001000000010000000001",
        88 => "0000000111100000000000111",
        
        96 => "0000000000000000100000001",  --- Instruccion de Subrutina
        97 => "0010000000000000000000001",
        98 => "0000000101000000000000001",
        99 => "0000000000000000100000001",
        100 => "0000010000000000000000001",
        101 => "0000000101000000000000001",
        102 => "0000000000000000100000001",
        103 => "0000001000000010000000001",
        104 => "0000000101000000000000001",
        105 => "0000000000001000000000001",
        106 => "0000000000000110100000001",
        107 => "0000000000000000010110001",
        108 => "0000000000001000000000001",
        109 => "0000000000000110100000001",
        110 => "0000000000000000010111001",
        111 => "0000000011100000000000011",

        112 => "0000000000000000100000001",  --- Instruccion de Retorno de Subrutina
        113 => "0010000000000000000000001",
        114 => "0000000000000110100000001",
        115 => "0000001000000000000000001",
        116 => "0000000000001000000000001",
        117 => "0000000000000110100000001",
        118 => "0000010000000000000000001",
        119 => "0000000000001000000000001",
        120 => "0000000011100000000000011",

        128 => "0000000000000000100000001",  --- Instruccion de Guardado de punteros
        129 => "0010000000000000000000001",
        130 => "0000000101000000000000001",
        131 => "0000000000000000100000001",
        132 => "0000010000000000000000001",
        133 => "0000000101000000000000001",
        134 => "0000000000000000100000001",
        135 => "0000001000000000000000001",
        136 => "0000000000000010100000001",
        137 => "0000000000000000011110001",
        138 => "0000000000000001000000001",
        139 => "0000000000000000011111001",
        140 => "0000000101000000000000011",

        144 => "0000000000000000100000001",  --- Instruccion de Carga de punteros Inmediata
        145 => "0010000000000000000000001",
        146 => "0000000101000000000000001",
        147 => "0000000000000000100000001",
        148 => "0000010000000000000000001",
        149 => "0000000101000000000000001",
        150 => "0000000000000000100000001",
        151 => "0000001000000000000000001",
        152 => "0000000101011000000000011",

        160 => "0000000000000000100000001",  --- Instruccion de Carga de punteros Directa
        161 => "0010000000000000000000001",
        162 => "0000000101000000000000001",
        163 => "0000000000000000100000001",
        164 => "0000010000000000000000001",
        165 => "0000000101000000000000001",
        166 => "0000000000000000100000001",
        167 => "0000001000000000000000001",
        168 => "0000000000000010100000001",
        169 => "0000010000000000000000001",
        170 => "0000000000000001000000001",
        171 => "0000001000000000000000001",
        172 => "0000000101011000000000011",

        176 => "0000000000000000100000001",  --- Instruccion de Guardado en pila de Acumulador
        177 => "0010000000000000000000001",
        178 => "0000000000001000000000001",
        179 => "0000000000000110100000001",
        180 => "0000000101000000011001111",

        192 => "0000000000000000100000001",  --- Instruccion de Guardado en pila de Punteros
        193 => "0010000000000000000000001",
        194 => "0000000000001000000000001",
        195 => "0000000000000110100000001",
        196 => "0000000000000000010010001",
        197 => "0000000000001000000000001",
        198 => "0000000000000110100000001",
        199 => "0000000000000000010011001",
        200 => "0000000101000000000000011",

        208 => "0000000000000000100000001",  --- Instruccion de Recuperado de pila Acumulador
        209 => "0010000000000000000000001",
        210 => "0000000000000110100000001",
        211 => "0000000101001000000000111",

        224 => "0000000000000000100000001",  --- Instruccion de Recuperado de pila Punteros
        225 => "0010000000000000000000001",
        226 => "0000000000000110100000001",
        227 => "0000001000000000000000001",
        228 => "0000000000001000000000001",
        229 => "0000000000000110100000001",
        230 => "0000010000000000000000001",
        231 => "0000000101010000000000001",
        232 => "0000000000001000000000011",

        240 => "0000000000000000100000001",  --- Instruccion de Salida de datos
        241 => "0010000000000000000000001",
        242 => "1000000101000000000000011",

        -- Finalizando a memoria com zeros
        others => "0000000000000000000000001"
    );

begin
    process(clk)
    begin
        if rising_edge(clk) then
            data <= mem(to_integer(unsigned(addr)));
        end if;
    end process;
end rtl;