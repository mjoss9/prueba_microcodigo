-- unidad secuencial de cálculo                        # S[0:30]  OK (USCE)

-- direccionamiento de memoria
-- inherente, inmediato, directo, indexado           # S[31:33] CC
-- [0,0,0] Secuencia de inicio
-- [0,0,1] Direccionamiento inherente
-- [0,1,0] Direccionamiento inmediato
-- [0,1,1] Direcciónamiento directo
-- [1,0,0] Direcciónamiento indexado

library ieee;
use ieee.std_logic_1164.all;

entity descodUSCE is
  port(
    in_s: in std_logic_vector(7 downto 0);
    out_s: out std_logic_vector(33 downto 0)
  );
end descodUSCE;
architecture arch of descodUSCE is
begin
  process(in_s) is
  begin
    case in_s is
      -- Instrucciones Logicas - Aritmeticas
        -- NEG
      when x"03" =>  out_s <= "0010010000000010000000011000010101"; -- neg A
      when x"13" =>  out_s <= "0010100000100010000000011000010101"; -- neg B
      when x"23" =>  out_s <= "0011000001000010000000011000010101"; -- neg C
      when x"33" =>  out_s <= "0110000010010010000000011000001011"; -- neg Mem
        -- NOT
      when x"04" =>  out_s <= "0010010000000010000000011000010100"; -- not A
      when x"14" =>  out_s <= "0010100000100010000000011000010100"; -- not B
      when x"24" =>  out_s <= "0011000001000010000000011000010100"; -- not C
      when x"34" =>  out_s <= "0110000010010010000000011000001010"; -- not Mem
        -- INC
      when x"43" =>  out_s <= "0010010000000011101000011000010001"; -- inc A
      when x"53" =>  out_s <= "0010100000100011101000011000010001"; -- inc B
      when x"63" =>  out_s <= "0011000001000011101000011000010001"; -- inc C
      when x"73" =>  out_s <= "0110000010010011101000011000001001"; -- inc Mem
        -- DEC
      when x"44" =>  out_s <= "0010010000000011101000011000010010"; -- dec A
      when x"54" =>  out_s <= "0010100000100011101000011000010010"; -- dec B
      when x"64" =>  out_s <= "0011000001000011101000011000010010"; -- dec C
      when x"74" =>  out_s <= "0110000010010011101000011000001100"; -- dec Mem 
        -- AND
      when x"55" =>  out_s <= "0010010110000010000000000000000000"; -- and AB
      when x"65" =>  out_s <= "0010011000000010000000000000000000"; -- and AC
      when x"95" =>  out_s <= "0010100100100010000000000000000000"; -- and BA
      when x"A5" =>  out_s <= "0010101000100010000000000000000000"; -- and BC
      when x"D5" =>  out_s <= "0011000101000010000000000000000000"; -- and CA
      when x"E5" =>  out_s <= "0011000111000010000000000000000000"; -- and CB
        -- OR
      when x"56" =>  out_s <= "0010010110000010000000001000000000"; -- or AB
      when x"66" =>  out_s <= "0010011000000010000000001000000000"; -- or AC
      when x"96" =>  out_s <= "0010100100100010000000001000000000"; -- or BA
      when x"A6" =>  out_s <= "0010101000100010000000001000000000"; -- or BC
      when x"D6" =>  out_s <= "0011000101000010000000001000000000"; -- or CA
      when x"E6" =>  out_s <= "0011000111000010000000001000000000"; -- or CB
        -- XOR
      when x"57" =>  out_s <= "0010010110000010000000010000000000"; -- xor AB
      when x"67" =>  out_s <= "0010011000000010000000010000000000"; -- xor AC
      when x"97" =>  out_s <= "0010100100100010000000010000000000"; -- xor BA
      when x"A7" =>  out_s <= "0010101000100010000000010000000000"; -- xor BC
      when x"D7" =>  out_s <= "0011000101000010000000010000000000"; -- xor CA
      when x"E7" =>  out_s <= "0011000111000010000000010000000000"; -- xor CB
        -- ADD
      when x"58" =>  out_s <= "0010010110000011101101011000011000"; -- add AB
      when x"68" =>  out_s <= "0010011000000011101101011000011000"; -- add AC
      when x"98" =>  out_s <= "0010100100100011101101011000011000"; -- add BA
      when x"A8" =>  out_s <= "0010101000100011101101011000011000"; -- add BC
      when x"D8" =>  out_s <= "0011000101000011101101011000011000"; -- add CA
      when x"E8" =>  out_s <= "0011000111000011101101011000011000"; -- add CB
        -- SUB
      when x"59" =>  out_s <= "0010010110000011101101011000011011"; -- sub AB
      when x"69" =>  out_s <= "0010011000000011101101011000011011"; -- sub AC
      when x"99" =>  out_s <= "0010100100100011101101011000011011"; -- sub BA
      when x"A9" =>  out_s <= "0010101000100011101101011000011011"; -- sub BC
      when x"D9" =>  out_s <= "0011000101000011101101011000011011"; -- sub CA
      when x"E9" =>  out_s <= "0011000111000011101101011000011011"; -- sub CB
        -- ADC
      when x"5A" =>  out_s <= "0010010110000011101101011000111000"; -- adc AB
      when x"6A" =>  out_s <= "0010011000000011101101011000111000"; -- adc AC
      when x"9A" =>  out_s <= "0010100100100011101101011000111000"; -- adc BA
      when x"AA" =>  out_s <= "0010101000100011101101011000111000"; -- adc BC
      when x"DA" =>  out_s <= "0011000101000011101101011000111000"; -- adc CA
      when x"EA" =>  out_s <= "0011000111000011101101011000111000"; -- adc CB
        -- SBC
      when x"5B" =>  out_s <= "0010010110000011101101011000111011"; -- sbc AB
      when x"6B" =>  out_s <= "0010011000000011101101011000111011"; -- sbc AC
      when x"9B" =>  out_s <= "0010100100100011101101011000111011"; -- sbc BA
      when x"AB" =>  out_s <= "0010101000100011101101011000111011"; -- sbc BC
      when x"DB" =>  out_s <= "0011000101000011101101011000111011"; -- sbc CA
      when x"EB" =>  out_s <= "0011000111000011101101011000111011"; -- sbc CB
        -- CMP
      when x"5C" =>  out_s <= "0010010110000011101101011000011011"; -- cmp AB
      when x"6C" =>  out_s <= "0010011000000011101101011000011011"; -- cmp AC
      when x"9C" =>  out_s <= "0010100100100011101101011000011011"; -- cmp BA
      when x"AC" =>  out_s <= "0010101000100011101101011000011011"; -- cmp BC
      when x"DC" =>  out_s <= "0011000101000011101101011000011011"; -- cmp CA
      when x"EC" =>  out_s <= "0011000111000011101101011000011011"; -- cmp CB
        -- Instrucciones con memoria
      when x"75" =>  out_s <= "0110010010000010000000000000000000"; -- and A_Mem
      when x"B5" =>  out_s <= "0110100010100010000000000000000000"; -- and B_Mem
      when x"F5" =>  out_s <= "0111000011000010000000000000000000"; -- and B_Mem

      when x"76" =>  out_s <= "0110010010000010000000001000000000"; -- or A_Mem
      when x"B6" =>  out_s <= "0110100010100010000000001000000000"; -- or B_Mem
      when x"F6" =>  out_s <= "0111000011000010000000001000000000"; -- or C_Mem

      when x"77" =>  out_s <= "0110010010000010000000010000000000"; -- xor A_Mem
      when x"B7" =>  out_s <= "0110100010100010000000010000000000"; -- xor B_Mem
      when x"F7" =>  out_s <= "0111000011000010000000010000000000"; -- xor C_Mem

      when x"78" =>  out_s <= "0110010010000011101101011000011000"; -- add A_Mem
      when x"B8" =>  out_s <= "0110100010100011101101011000011000"; -- add B_Mem
      when x"F8" =>  out_s <= "0111000011000011101101011000011000"; -- add C_Mem

      when x"79" =>  out_s <= "0110010010000011101101011000011011"; -- sub A_Mem
      when x"B9" =>  out_s <= "0110100010100011101101011000011011"; -- sub B_Mem
      when x"F9" =>  out_s <= "0111000011000011101101011000011011"; -- sub C_Mem

      when x"7A" =>  out_s <= "0110010010000011101101011000111000"; -- adc A_Mem
      when x"BA" =>  out_s <= "0110100010100011101101011000111000"; -- adc B_Mem
      when x"FA" =>  out_s <= "0111000011000011101101011000111000"; -- adc C_Mem

      when x"7B" =>  out_s <= "0110010010000011101101011000111011"; -- sbc A_Mem
      when x"BB" =>  out_s <= "0110100010100011101101011000111011"; -- sbc B_Mem
      when x"FB" =>  out_s <= "0111000011000011101101011000111011"; -- sbc C_Mem

      when x"7C" =>  out_s <= "0110010010000011101101011000011011"; -- cmp A_Mem
      when x"BC" =>  out_s <= "0110100010100011101101011000011011"; -- cmp B_Mem
      when x"FC" =>  out_s <= "0111000011000011101101011000011011"; -- cmp C_Mem

      -- Instrucciones Control
      when x"00" =>  out_s <= "0000000000000000000000011000010000"; -- nop
      when x"20" =>  out_s <= "0010000000000000000100011000010000"; -- clc
      when x"30" =>  out_s <= "0010000000000000000110011000010000"; -- clv
      when x"90" =>  out_s <= "0010000000000000100000011000010000"; -- sec
      when x"A0" =>  out_s <= "0010000000000000110000011000010000"; -- sev

        -- Instrucciones de limpieza de datos
      when x"01" =>  out_s <= "0010010000000010000000011000000000"; -- clr A
      when x"11" =>  out_s <= "0010100000100010000000011000000000"; -- clr B
      when x"21" =>  out_s <= "0011000001000010000000011000000000"; -- clr C
          -- Instrucciones de limpieza de datos en memoria
      when x"31" =>  out_s <= "0110000000010010000000011000000000"; -- clr Mem
      
      -- Instrucciones Entrada de datos
      when x"02" =>  out_s <= "0010010000000010000000011000001000"; -- in A
      when x"12" =>  out_s <= "0010100000000010000000011000001000"; -- in B
      when x"22" =>  out_s <= "0011000000000010000000011000001000"; -- in C
        -- Instrucciones de carga de memoria
      when x"71" =>  out_s <= "0110010010000010000000011000001000"; -- lda A_Mem
      when x"B1" =>  out_s <= "0110100010000010000000011000001000"; -- lda A_Mem
      when x"F1" =>  out_s <= "0111000010000010000000011000001000"; -- lda A_Mem
        -- Instrucciones de guardado en memoria
      when x"72" =>  out_s <= "0110000000010000000000011000010000"; -- sta A_Mem
      when x"B2" =>  out_s <= "0110000000110000000000011000010000"; -- sta B_Mem
      when x"F2" =>  out_s <= "0110000001010000000000011000010000"; -- sta C_Mem

      -- Instrucciones Rotamiento - Desplazamiento
        -- Rotaciones
      when x"0D" =>  out_s <= "0010010000000010000101100000010000"; -- rod A
      when x"0E" =>  out_s <= "0010010000000010000101100010010000"; -- roi A
      when x"4D" =>  out_s <= "0010010000000010000101100001010000"; -- rcd A
      when x"4E" =>  out_s <= "0010010000000010000101100011010000"; -- rci A

      when x"1D" =>  out_s <= "0010100000100010000101100000010000"; -- rod B
      when x"1E" =>  out_s <= "0010100000100010000101100010010000"; -- roi B
      when x"5D" =>  out_s <= "0010100000100010000101100001010000"; -- rcd B
      when x"5E" =>  out_s <= "0010100000100010000101100011010000"; -- rci B

      when x"2D" =>  out_s <= "0011000001000010000101100000010000"; -- rod C
      when x"2E" =>  out_s <= "0011000001000010000101100010010000"; -- roi C
      when x"6D" =>  out_s <= "0011000001000010000101100001010000"; -- rcd C
      when x"6E" =>  out_s <= "0011000001000010000101100011010000"; -- rci C
          -- Rotaciones con memoria
      when x"3D" =>  out_s <= "0110000010010010000101100000001000"; -- rod Mem
      when x"3E" =>  out_s <= "0110000010010010000101100010001000"; -- roi Mem
      when x"7D" =>  out_s <= "0110000010010010000101100001001000"; -- rcd Mem
      when x"7E" =>  out_s <= "0110000010010010000101100011001000"; -- rci Mem

        -- Desplazamientos
      when x"8D" =>  out_s <= "0010010000000010000101100100010000"; -- dad A
      when x"8E" =>  out_s <= "0010010000000010000101100110010000"; -- dai A
      when x"CD" =>  out_s <= "0010010000000010000101100101010000"; -- dld A

      when x"9D" =>  out_s <= "0010100000100010000101100100010000"; -- dad B
      when x"9E" =>  out_s <= "0010100000100010000101100110010000"; -- dai B
      when x"DD" =>  out_s <= "0010100000100010000101100101010000"; -- dld B

      when x"AD" =>  out_s <= "0011000001000010000101100100010000"; -- dad C
      when x"AE" =>  out_s <= "0011000001000010000101100110010000"; -- dai C
      when x"ED" =>  out_s <= "0011000001000010000101100101010000"; -- dld C
          -- Desplazamientos con memoria
      when x"BD" =>  out_s <= "0110000010010010000101100100001000"; -- dad Mem
      when x"BE" =>  out_s <= "0110000010010010000101100110001000"; -- dai Mem
      when x"FD" =>  out_s <= "0110000010010010000101100101001000"; -- dld Mem

        -- Trasferencias
      when x"91" =>  out_s <= "0010100000000010000000011000001000"; -- lda BA
      when x"D1" =>  out_s <= "0011000000000010000000011000001000"; -- lda CA
      when x"51" =>  out_s <= "0010010000100010000000011000001000"; -- lda AB
      when x"E1" =>  out_s <= "0011000000100010000000011000001000"; -- lda CB
      when x"61" =>  out_s <= "0010010001000010000000011000001000"; -- lda AC
      when x"A1" =>  out_s <= "0010100001000010000000011000001000"; -- lda BC

      when others => out_s <= "0000000000000000000000000000000000";
    end case;
  end process;
end arch;